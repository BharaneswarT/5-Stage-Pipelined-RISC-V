module imm_gen(
	input [31:0] instr,
	input [7:0] opcode,
	output reg [31:0] imm
	);
	
	always @(*) begin
        case(opcode)
            // I-type instruction (loads, jalr, immediate arith)
            7'b0000011, 7'b0010011, 7'b1100111: imm = {{20{instr[31]}}, instr[31:20]};
            
            // S-type instruction(stores)
            7'b0100011: imm = {{20{instr[31]}}, instr[31:25], instr[11:7]};
            
            // B-type instr(branches)
            7'b1100011: imm = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
            
            // U-type instr (lui/auipc)
            7'b0110111, 7'b0010111: imm = {instr[31:12], 12'b0};
            
            // J-type instr(jal)
            7'b1101111: imm = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
            
            default: imm = 0;  // R-type instr
            
        endcase
    end
endmodule
